module Mux4to1 (
    input [7:0] D0, D1, D2, D3,
    input [1:0] Addr,
    output reg [7:0] Q
);

always @(*) begin 
    case (Addr)
        2'b00: Q = D0;
        2'b01: Q = D1;
        2'b10: Q = D2;
        2'b11: Q = D3;
        default: Q = 8'b00000000;
    endcase
end

endmodule
